library verilog;
use verilog.vl_types.all;
entity perity_check_vlg_vec_tst is
end perity_check_vlg_vec_tst;
