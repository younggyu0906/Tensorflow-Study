library verilog;
use verilog.vl_types.all;
entity hw2logic_vlg_vec_tst is
end hw2logic_vlg_vec_tst;
