library verilog;
use verilog.vl_types.all;
entity comparator_vlg_vec_tst is
end comparator_vlg_vec_tst;
