library verilog;
use verilog.vl_types.all;
entity ringCount_vlg_vec_tst is
end ringCount_vlg_vec_tst;
