library verilog;
use verilog.vl_types.all;
entity parity_vlg_vec_tst is
end parity_vlg_vec_tst;
