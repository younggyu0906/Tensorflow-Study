library verilog;
use verilog.vl_types.all;
entity add4_vlg_vec_tst is
end add4_vlg_vec_tst;
