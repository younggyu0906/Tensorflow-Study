library verilog;
use verilog.vl_types.all;
entity reg_combin_vlg_vec_tst is
end reg_combin_vlg_vec_tst;
