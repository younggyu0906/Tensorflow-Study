library verilog;
use verilog.vl_types.all;
entity combosys_vlg_check_tst is
    port(
        o1              : in     vl_logic;
        o2              : in     vl_logic;
        o3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end combosys_vlg_check_tst;
