library verilog;
use verilog.vl_types.all;
entity or2test_vlg_vec_tst is
end or2test_vlg_vec_tst;
