library verilog;
use verilog.vl_types.all;
entity ex02_vlg_vec_tst is
end ex02_vlg_vec_tst;
