library verilog;
use verilog.vl_types.all;
entity signal_lamp_vlg_vec_tst is
end signal_lamp_vlg_vec_tst;
