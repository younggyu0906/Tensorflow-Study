library verilog;
use verilog.vl_types.all;
entity claDesign_vlg_vec_tst is
end claDesign_vlg_vec_tst;
