library verilog;
use verilog.vl_types.all;
entity system_vlg_vec_tst is
end system_vlg_vec_tst;
