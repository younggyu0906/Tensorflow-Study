library verilog;
use verilog.vl_types.all;
entity kygmin1_vlg_vec_tst is
end kygmin1_vlg_vec_tst;
