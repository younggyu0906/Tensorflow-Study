library verilog;
use verilog.vl_types.all;
entity laundry_vlg_vec_tst is
end laundry_vlg_vec_tst;
