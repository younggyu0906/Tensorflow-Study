library verilog;
use verilog.vl_types.all;
entity signal_lamp_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end signal_lamp_vlg_sample_tst;
