library verilog;
use verilog.vl_types.all;
entity sys_var_vlg_vec_tst is
end sys_var_vlg_vec_tst;
