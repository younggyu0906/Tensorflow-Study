library verilog;
use verilog.vl_types.all;
entity and3input_vlg_check_tst is
    port(
        o               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end and3input_vlg_check_tst;
