library verilog;
use verilog.vl_types.all;
entity cla4_vlg_vec_tst is
end cla4_vlg_vec_tst;
