library verilog;
use verilog.vl_types.all;
entity nor4test_vlg_vec_tst is
end nor4test_vlg_vec_tst;
