library verilog;
use verilog.vl_types.all;
entity andlogic_vlg_vec_tst is
end andlogic_vlg_vec_tst;
