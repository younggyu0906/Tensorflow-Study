library verilog;
use verilog.vl_types.all;
entity jk_counter2_vlg_vec_tst is
end jk_counter2_vlg_vec_tst;
