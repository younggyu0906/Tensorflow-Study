library verilog;
use verilog.vl_types.all;
entity hw02_vlg_check_tst is
    port(
        agtb            : in     vl_logic;
        altb            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hw02_vlg_check_tst;
