library verilog;
use verilog.vl_types.all;
entity bcdAdder_vlg_vec_tst is
end bcdAdder_vlg_vec_tst;
