library verilog;
use verilog.vl_types.all;
entity hw02_vlg_vec_tst is
end hw02_vlg_vec_tst;
