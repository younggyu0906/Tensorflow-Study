library verilog;
use verilog.vl_types.all;
entity decoder24_vlg_vec_tst is
end decoder24_vlg_vec_tst;
