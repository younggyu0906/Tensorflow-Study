library verilog;
use verilog.vl_types.all;
entity hw3decoder24_vlg_vec_tst is
end hw3decoder24_vlg_vec_tst;
