library verilog;
use verilog.vl_types.all;
entity or2test_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end or2test_vlg_check_tst;
