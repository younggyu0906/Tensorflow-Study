library verilog;
use verilog.vl_types.all;
entity comp_vlg_check_tst is
    port(
        equal           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end comp_vlg_check_tst;
