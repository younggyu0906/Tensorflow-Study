library verilog;
use verilog.vl_types.all;
entity and2test_vlg_vec_tst is
end and2test_vlg_vec_tst;
