library verilog;
use verilog.vl_types.all;
entity logic_vlg_vec_tst is
end logic_vlg_vec_tst;
