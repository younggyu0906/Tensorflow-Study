library verilog;
use verilog.vl_types.all;
entity system_vlg_check_tst is
    port(
        y_out           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end system_vlg_check_tst;
