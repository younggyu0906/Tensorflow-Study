library verilog;
use verilog.vl_types.all;
entity jk_counter_vlg_vec_tst is
end jk_counter_vlg_vec_tst;
