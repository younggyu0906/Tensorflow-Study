library verilog;
use verilog.vl_types.all;
entity and3input_vlg_vec_tst is
end and3input_vlg_vec_tst;
