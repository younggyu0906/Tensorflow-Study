library verilog;
use verilog.vl_types.all;
entity sys_var_vlg_check_tst is
    port(
        l               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sys_var_vlg_check_tst;
