library verilog;
use verilog.vl_types.all;
entity nor_sys_vlg_check_tst is
    port(
        c               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end nor_sys_vlg_check_tst;
