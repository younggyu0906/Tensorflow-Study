library verilog;
use verilog.vl_types.all;
entity KYGLJY_Robot_vlg_vec_tst is
end KYGLJY_Robot_vlg_vec_tst;
