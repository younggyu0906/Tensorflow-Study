library verilog;
use verilog.vl_types.all;
entity logic2_vlg_check_tst is
    port(
        y_out           : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end logic2_vlg_check_tst;
