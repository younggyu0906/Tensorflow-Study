library verilog;
use verilog.vl_types.all;
entity kygmaxmin2_vlg_vec_tst is
end kygmaxmin2_vlg_vec_tst;
