library verilog;
use verilog.vl_types.all;
entity kygmin2 is
    port(
        a               : in     vl_logic_vector(7 downto 0);
        b               : in     vl_logic_vector(7 downto 0);
        y_out           : out    vl_logic_vector(7 downto 0)
    );
end kygmin2;
