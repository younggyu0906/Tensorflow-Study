library verilog;
use verilog.vl_types.all;
entity kygmaxmin_vlg_vec_tst is
end kygmaxmin_vlg_vec_tst;
