library verilog;
use verilog.vl_types.all;
entity apollo_vlg_vec_tst is
end apollo_vlg_vec_tst;
