library verilog;
use verilog.vl_types.all;
entity nor_sys_vlg_vec_tst is
end nor_sys_vlg_vec_tst;
