library verilog;
use verilog.vl_types.all;
entity combosys_vlg_vec_tst is
end combosys_vlg_vec_tst;
