library verilog;
use verilog.vl_types.all;
entity logic2_vlg_vec_tst is
end logic2_vlg_vec_tst;
