library verilog;
use verilog.vl_types.all;
entity adder_16_vlg_vec_tst is
end adder_16_vlg_vec_tst;
