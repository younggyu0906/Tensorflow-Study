library verilog;
use verilog.vl_types.all;
entity reg_decom_vlg_vec_tst is
end reg_decom_vlg_vec_tst;
