library verilog;
use verilog.vl_types.all;
entity hw01_vlg_check_tst is
    port(
        agtb            : in     vl_logic;
        altb            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end hw01_vlg_check_tst;
