library verilog;
use verilog.vl_types.all;
entity jk_flipflop_vlg_vec_tst is
end jk_flipflop_vlg_vec_tst;
