library verilog;
use verilog.vl_types.all;
entity hw01_vlg_vec_tst is
end hw01_vlg_vec_tst;
