library verilog;
use verilog.vl_types.all;
entity kygmin2_vlg_vec_tst is
end kygmin2_vlg_vec_tst;
