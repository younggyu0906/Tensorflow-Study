library verilog;
use verilog.vl_types.all;
entity rcaAdder_vlg_vec_tst is
end rcaAdder_vlg_vec_tst;
