library verilog;
use verilog.vl_types.all;
entity kygmaxmin3_vlg_vec_tst is
end kygmaxmin3_vlg_vec_tst;
