library verilog;
use verilog.vl_types.all;
entity reg4_vlg_vec_tst is
end reg4_vlg_vec_tst;
